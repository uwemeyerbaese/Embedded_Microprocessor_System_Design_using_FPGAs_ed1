-- ------------------------------------------------
-- VHDL STD 1076-1993 keywords
-- ------------------------------------------------
ABS
ACCESS
AFTER
ALIAS
ALL
AND
ARCHITECTURE
ARRAY
ASSERT
ATTRIBUTE

BEGIN
BLOCK
BODY
BUFFER
BUS

CASE
COMPONENT
CONFIGURATION
CONSTANT

DISCONNECT
DOWNTO

ELSE
ELSIF
END
ENTITY
EXIT

FILE
FOR
FUNCTION

GENERATE
GENERIC
GROUP
GUARDED

IF
IMPURE
IN
INERTIAL
INOUT
IS

LABEL
LIBRARY
LINKAGE
LITERAL
LOOP

MAP
MOD

NAND
NEW
NEXT
NOR
NOT
NULL

OF
ON
OPEN
OR
OTHERS
OUT

PACKAGE
PORT
POSTPONED
PROCEDURE
PROCESS
PURE

RANGE
RECORD
REGISTER
REJECT
REM
REPORT
RETURN
ROL
ROR

SELECT
SEVERITY
SHARED
SIGNAL
SLA
SLL
SRA
SRL
SUBTYPE

THEN
TO
TRANSPORT
TYPE

UNAFFECTED
UNITS
UNTIL
USE

VARIABLE

WAIT
WHEN
WHILE
WITH

XNOR
XOR
