// ------------------------------------------------
// Verilog STD 1364-1995 keywords
// ------------------------------------------------

always
and
assign

begin
buf
bufif0
bufif1

case
casex
casez
cmos

deassign
default
defparam
disable

edge
else
end
endcase
endmodule
endfunction
endprimitive
endspecify
endtable
endtask
event

for
force
forever
fork
function

highz0
highz1

if
ifnone
initial
inout
input
integer

join

large

macromodule
medium
module

nand
negedge
nmos
nor
not
notif0
notif1

or
output

parameter
pmos
posedge
primitive
pull0
pull1
pullup
pulldown

rcmos
real
realtime
reg
release
repeat
rnmos
rpmos
rtran
rtranif0
rtranif1

scalared
small
specify
specparam
strong0
strong1
supply0
supply1

table
task
time
tran
tranif0
tranif1
tri
tri0
tri1
triand
trior
trireg

vectored

wait
wand
weak0
weak1
while
wire
wor

xnor
xor
