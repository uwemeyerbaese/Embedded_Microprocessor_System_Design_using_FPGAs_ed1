-- ------------------------------------------------
-- VHDL STD 1076-2008 keywords
-- ------------------------------------------------
ABS
ACCESS
AFTER
ALIAS
ALL
AND
ARCHITECTURE
ARRAY
ASSERT
ASSUME
ASSUME_GUARANTEE
ATTRIBUTE

BEGIN
BLOCK
BODY
BUFFER
BUS

CASE
COMPONENT
CONFIGURATION
CONSTANT
CONTEXT
COVER

DEFAULT
DISCONNECT
DOWNTO

ELSE
ELSIF
END
ENTITY
EXIT

FAIRNESS
FILE
FOR
FORCE
FUNCTION

GENERATE
GENERIC
GROUP
GUARDED

IF
IMPURE
IN
INERTIAL
INOUT
IS

LABEL
LIBRARY
LINKAGE
LITERAL
LOOP

MAP
MOD

NAND
NEW
NEXT
NOR
NOT
NULL

OF
ON
OPEN
OR
OTHERS
OUT

PACKAGE
PARAMETER
PORT
POSTPONED
PROCEDURE
PROCESS
PROPERTY
PROTECTED
PURE

RANGE
RECORD
REGISTER
REJECT
RELEASE
REM
REPORT
RESTRICT
RESTRICT_GUARANTEE
RETURN
ROL
ROR

SELECT
SEQUENCE
SEVERITY
SHARED
SIGNAL
SLA
SLL
SRA
SRL
STRONG
SUBTYPE

THEN
TO
TRANSPORT
TYPE

UNAFFECTED
UNITS
UNTIL
USE

VARIABLE
VMODE
VPROP
VUNIT

WAIT
WHEN
WHILE
WITH

XNOR
XOR
